//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW2AR-LV18QN88PC8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Wed Jul 24 02:35:37 2024

module rom_font_1bit (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [13:0] ad;

wire [30:0] prom_inst_0_dout_w;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h00081C3E7F7F7F367EFFE7C3FFDBFF7E7E8199BD81A5817E0000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000183C3C1800003E1C3E7F3E1C08083E1C3E7F7F1C3E1C00081C3E7F3E1C08;
defparam prom_inst_0.INIT_RAM_02 = 256'h1E333333BEF0E0F0FFC399BDBD99C3FF003C664242663C00FFFFE7C3C3E7FFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'h995A3CE7E73C5A990367E6C6C6FEC6FE070F0E0C0CFCCCFC187E183C6666663C;
defparam prom_inst_0.INIT_RAM_04 = 256'h0066006666666666183C7E18187E3C180040707C7F7C70400001071F7F1F0701;
defparam prom_inst_0.INIT_RAM_05 = 256'hFF183C7E187E3C18007E7E7E000000001E331C36361CC67C00D8D8D8DEDBDBFE;
defparam prom_inst_0.INIT_RAM_06 = 256'h00000C067F060C00000018307F30180000183C7E1818181800181818187E3C18;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000183C7EFFFF000000FFFF7E3C180000002466FF66240000007F0303030000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0036367F367F36360000000000363636000C000C0C1E1E0C0000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000030606006E333B6E1C361C0063660C18336300000C1F301E033E0C;
defparam prom_inst_0.INIT_RAM_0A = 256'h00000C0C3F0C0C000000663CFF3C660000060C1818180C0600180C0606060C18;
defparam prom_inst_0.INIT_RAM_0B = 256'h000103060C183060000C0C0000000000000000003F000000060C0C0000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h001E33301C30331E003F33061C30331E003F0C0C0C0C0E0C003E676F7B73633E;
defparam prom_inst_0.INIT_RAM_0D = 256'h000C0C0C1830333F001E33331F03061C001E3330301F033F0078307F33363C38;
defparam prom_inst_0.INIT_RAM_0E = 256'h060C0C00000C0C00000C0C00000C0C00000E18303E33331E001E33331E33331E;
defparam prom_inst_0.INIT_RAM_0F = 256'h000C000C1830331E00060C1830180C0600003F00003F000000180C0603060C18;
defparam prom_inst_0.INIT_RAM_10 = 256'h003C66030303663C003F66663E66663F0033333F33331E0C001E037B7B7B633E;
defparam prom_inst_0.INIT_RAM_11 = 256'h007C66730303663C000F06161E16467F007F46161E16467F001F36666666361F;
defparam prom_inst_0.INIT_RAM_12 = 256'h006766361E366667001E333330303078001E0C0C0C0C0C1E003333333F333333;
defparam prom_inst_0.INIT_RAM_13 = 256'h001C36636363361C006363737B6F67630063636B7F7F7763007F66460606060F;
defparam prom_inst_0.INIT_RAM_14 = 256'h001E33380E07331E006766363E66663F00381E3B3333331E000F06063E66663F;
defparam prom_inst_0.INIT_RAM_15 = 256'h0063777F6B636363000C1E3333333333003F333333333333001E0C0C0C0C2D3F;
defparam prom_inst_0.INIT_RAM_16 = 256'h001E06060606061E007F664C1831637F001E0C0C1E3333330063361C1C366363;
defparam prom_inst_0.INIT_RAM_17 = 256'hFF000000000000000000000063361C08001E18181818181E00406030180C0603;
defparam prom_inst_0.INIT_RAM_18 = 256'h001E3303331E0000003B66663E060607006E333E301E00000000000000180C0C;
defparam prom_inst_0.INIT_RAM_19 = 256'h1F303E33336E0000000F06060F06361C001E033F331E0000006E33333E303038;
defparam prom_inst_0.INIT_RAM_1A = 256'h0067361E366606071E33333030300030001E0C0C0C0E000C006766666E360607;
defparam prom_inst_0.INIT_RAM_1B = 256'h001E3333331E000000333333331F000000636B7F7F330000001E0C0C0C0C0C0E;
defparam prom_inst_0.INIT_RAM_1C = 256'h001F301E033E0000000F06666E3B000078303E33336E00000F063E66663B0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h00367F7F6B630000000C1E3333330000006E33333333000000182C0C0C3E0C08;
defparam prom_inst_0.INIT_RAM_1E = 256'h00380C0C070C0C38003F260C193F00001F303E33333300000063361C36630000;
defparam prom_inst_0.INIT_RAM_1F = 256'h007F6363361C08000000000000003B6E00070C0C380C0C070018181800181818;
defparam prom_inst_0.INIT_RAM_20 = 256'h00FC667C603CC37E001E033F331E0038007E3333330033001E30181E3303331E;
defparam prom_inst_0.INIT_RAM_21 = 256'h1C301E03031E0000007E333E301E0C0C007E333E301E0007007E333E301E0033;
defparam prom_inst_0.INIT_RAM_22 = 256'h001E0C0C0C0E0033001E033F331E0007001E033F331E0033003C067E663CC37E;
defparam prom_inst_0.INIT_RAM_23 = 256'h00333F331E000C0C0063637F63361C63001E0C0C0C0E0007003C1818181C633E;
defparam prom_inst_0.INIT_RAM_24 = 256'h001E33331E00331E007333337F33367C00FE33FE30FE0000003F061E063F0038;
defparam prom_inst_0.INIT_RAM_25 = 256'h007E333333000700007E33333300331E001E33331E000700001E33331E003300;
defparam prom_inst_0.INIT_RAM_26 = 256'h18187E03037E1818001E33333333003300183C66663C18C31F303E3333003300;
defparam prom_inst_0.INIT_RAM_27 = 256'h0E1B18183C18D870E363F3635F33331F0C0C3F0C3F1E3333003F67060F26361C;
defparam prom_inst_0.INIT_RAM_28 = 256'h007E333333003800001E33331E003800001E0C0C0C0E001C007E333E301E0038;
defparam prom_inst_0.INIT_RAM_29 = 256'h00003E001C36361C00007E007C36363C00333B3F3733003F003333331F001F00;
defparam prom_inst_0.INIT_RAM_2A = 256'hF03366CC7B3363C3000030303F000000000003033F000000001E3303060C000C;
defparam prom_inst_0.INIT_RAM_2B = 256'h00003366CC6633000000CC663366CC000018181818001818C0F3F6ECDB3363C3;
defparam prom_inst_0.INIT_RAM_2C = 256'h181818181818181877DBEEDB77DBEEDB55AA55AA55AA55AA1144114411441144;
defparam prom_inst_0.INIT_RAM_2D = 256'h6C6C6C7F000000006C6C6C6F6C6C6C6C1818181F181F18181818181F18181818;
defparam prom_inst_0.INIT_RAM_2E = 256'h6C6C6C6F607F00006C6C6C6C6C6C6C6C6C6C6C6F606F6C6C1818181F181F0000;
defparam prom_inst_0.INIT_RAM_2F = 256'h1818181F000000000000001F181F18180000007F6C6C6C6C0000007F606F6C6C;
defparam prom_inst_0.INIT_RAM_30 = 256'h181818F818181818181818FF00000000000000FF18181818000000F818181818;
defparam prom_inst_0.INIT_RAM_31 = 256'h6C6C6CEC6C6C6C6C181818F818F81818181818FF18181818000000FF00000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h6C6C6CEF00FF0000000000FF00EF6C6C6C6C6CEC0CFC0000000000FC0CEC6C6C;
defparam prom_inst_0.INIT_RAM_33 = 256'h000000FF00FF18186C6C6CEF00EF6C6C000000FF00FF00006C6C6CEC0CEC6C6C;
defparam prom_inst_0.INIT_RAM_34 = 256'h000000FC6C6C6C6C6C6C6CFF00000000181818FF00FF0000000000FF6C6C6C6C;
defparam prom_inst_0.INIT_RAM_35 = 256'h6C6C6CFF6C6C6C6C6C6C6CFC00000000181818F818F80000000000F818F81818;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF181818F8000000000000001F18181818181818FF18FF1818;
defparam prom_inst_0.INIT_RAM_37 = 256'h00000000FFFFFFFFF0F0F0F0F0F0F0F00F0F0F0F0F0F0F0FFFFFFFFF00000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0036363636367F000003030303333F0003031F331F331E00006E3B133B6E0000;
defparam prom_inst_0.INIT_RAM_39 = 256'h00181818183B6E0003063E6666666600000E1B1B1B7E0000003F33060C06333F;
defparam prom_inst_0.INIT_RAM_3A = 256'h001E33333E180C38007736366363361C001C36637F63361C3F0C1E33331E0C3F;
defparam prom_inst_0.INIT_RAM_3B = 256'h003333333333331E001C06031F03061C03067EDBDB7E306000007EDBDB7E0000;
defparam prom_inst_0.INIT_RAM_3C = 256'h003F00180C060C18003F00060C180C06003F000C0C3F0C0C00003F003F003F00;
defparam prom_inst_0.INIT_RAM_3D = 256'h00003B6E003B6E00000C0C003F000C0C0E1B1B18181818181818181818D8D870;
defparam prom_inst_0.INIT_RAM_3E = 256'h383C3637303030F000000018000000000000001818000000000000001C36361C;
defparam prom_inst_0.INIT_RAM_3F = 256'h000000000000000000003C3C3C3C00000000001E060C180E000000363636361E;

endmodule //rom_font_1bit
